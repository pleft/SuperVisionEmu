                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           H�Z� �h ��n ��m � �k ���i �i ��k �  m��i �r� ���i ��d�l ���j �i �i ��k � � �h ��m  m��j �j �j ��l � ��m ��h  m��j �D� ���� �� ���i ���m �k � � �h  ���k i�k �  m��l � ��h  ���l 8��l �  m��l �T� ����z�hL� ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<3<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                        ��      �*V�V�V�V�V���*      �?�?      H��!��"�(� �)� C�h`Hڭt������ ���(i�&0�&��( Y���� � J�����h`Hڭ@�,���@� ���A�i
�I���Y�2��a�����h`	
H�Z�
�8�@���1�l�琍b� �`�,@���b���@�@�u� z� T���
z�h`HZ�! �Q��A��I�u�Y�u�2��azh`H��"��-��#��
 t��5 4��0 ��+��#�#� l�� �����#��
 <�� �� ˃h`H8��"��8�#����	P��! �� �! ���! h`H��! h`H8��"�8�#����	P��! ���! ���! h`H��! h`H8�"��8��#���	P�	�! ���! ��
�! h`H��! h`H8��"�8��#���	P��! ���! ���! h`H�Z�@�?� �`�,@�+�a�& � A� ����� �`�,@��
�( Y�2��a���� Y�z�h`HZ�A� �I��Y�i��!�v��" h�����  L�zh`HZ�A� �I��Y�i��!�v��" �� C�zh`H�Y� Q�� ��h`HZ�Q
���$ ȹ�% � �$}A0�&�A��$}Iɀ�	� ��I� ��zh`�h�-@�@`HZ�Y�Ay��0�&��A���}I� �	ɀ��I� ��zh`HZ A�(���$zh`HZ�
�����$ ȹ���% �� �$ȑ$zh`H�Z B��"JJJ����!J� څ��
�������������z�h`H� J��JJJ�h`H�
� �


�h`HZ B��"JJJ����!J� Ʌ��
�������������zh`H� ��
 �!�� �
8�!� �!�
�( h�h`H�Z� �. �!�6 �"�> �';� �F � ���l�0�. �!�6 �"�> � � � ��� �	��ж� ��z�h`Hڮ �. �!�6 �"�> � �F � e�� � e�� �	���Ӣ ���h`H� ��
 �!�� �
8�!� �! ��h` B� A���
�2�1� ˇ��# �`� A���
��1� ˇ��# �`� �& `���& `�Z8�2���8�2��g ����i����� � ���0�r  �Žh�-����& z�`H�Z�#��� ���	� �L���
�L������g ���	��i���ƚ���j�ƚ����P�s ���&L������P�s ��ɯ��P�s ���}��P�s ���d���s �d�d�2����P������r ��0�r  �� �� �� �����& z�h`���8�
��h�-# �# �i
�`�h�-���`��!��" C� �� �� ��`HZ�&�����!��"�?� � ��� Lݩ *� �`�,v������v�v� �w��}���zh`Hڭv�"� �`�,v���� w��h�-v�v�����h`H�w� �}���!��" C�h`�	�!� �"�B�  Lݩ *� �`HZ�l
��ˑ�$ ȹˑ�% �n�$�c��n�?�� � ��zh`HZ�l
��ۑ�$ ȹۑ�% �n
��$� ȱ$� �o�� ��c��o�n� #��ozh`HZ G��! �2� w��" �?zh` ���" �?zh`�l
��
��$ ȹ
��% �" �$`�l
����$ ȹ��% �?�$`������# ��� �` P�`H�t����l���0�+����� ���#�h`HZ�����.�l
�����$ ȹ���% �" �$�c��!  ���" ��" ���+zh`H�Z� �`�,�����J������l
����� ��$ ȹ��� ��% �" �$������ �����! ���! �
���z�h`H�Z� �`�,���������� ���! �
���� ��z�h`H�Z� �`�,# ������# �# �i
� ���! �
���� ��z�h`H�! �� �LO��� ��LO��� K�LO��� Q�LO��� K�LO��� ��LO��� K�LO��� ��LO�� � K�LO��!� K�LO��"� ��LO��#� ��LO��'� K�LO� _����'��� ���! ��h`H�! ���'��� _���� z��! ��h`H�! �� _������� ��h`HZ�! �� _����iJ��� A��
����� U�����j� �� �zh`H�Z���3� �`�,��"��� �� _��`�,���( Kϼ��
�������z�h`H�Z�# �G� �`�,# �6�i
����' �� _��8�
��`�,# ��i
��( Kϼ��
����8�
���耻z�h`H���� ��L)��� ��L)��� ��L)��� /�L)��� /�L)��� ��L)��� ��L)��� z�L)��	� ��L)��
� ��L)��� ��L)��� ��L)��� +�L)��� +�L)��� +�L)��� ��L)��� "�L)��� g�L)��� ��L)��� ��L)��� =�L)��� =�L)��� h�L)��� h�L)��� ��L)��� ��L)��� ��L)��� V�L)��� V�L)��� V�L)��� V�L)�� � ��L)��!� ��L)��"� ��L)��#� ��L)��$� �L)��%� F�L)��&� ��L)��'� �րA�(� ��L)��)� ��L)��*� ��L)��+� �L)��,� �Ԁ�-� �׀�.� �h`]�j�v��������������������ɏԏߏ} � � ���	��.�:�PRESSaSTARTa$PRESSaSTART$CONTINUE$END$BEAM$SCORE$NUM$READY$GAMEaaOVER$PAUSE$STAGEaONE$STAGEaTWO$STAGEaTHREE$STAGEaFOUR$STAGEaFIVE$STAGEaSIX$ENTERaYOURaNAME$CHOOSEaaMISSION$CONGRATULATIONaYOU$SEEaYOUaNEXTaTIME$HIGHaSCOREa$YOURaSCOREa$������$�ĝ����+�1�q����1�9�y�����9�]�e�u������)�A�����¢ڢ�
�$�<�L������������0�Y�u���ƥ��#�d���(�����`�Ȩب����� �@�P�`����������x�|��p�3�������󲧳%�6�V�f���V���6�đ

	
8' CDEFGHIJKLMN	
	
	
	

	c   c	
		
		
	c     ccc  c������(�@�@�D�f�������Ԓ��	
c	
cc	
c	
c	
 !#cc*�/�2�5�8�;�?�B�D�G�I�K�P�S�V�Y�`���������Ɠ˓Γדړޓ���H�M�Q�U�Y�\�a�d�h�m�q�w�{������������"�*�1�7�H�M�T�Y�_����&�,�2�4�>�B�F�L�P�U�Ӗؖܖ������������	�����"�%�*�/�3�;�;�?�F�Q�b����f�W�T��������͔��������ccccccccccc
cccc
cc$PV\06<ZPJBLZR( PH<4FP$X(2	cc
cc	cccccccccPHX<^4Z((RFFZ(<<F0\(ZPPZ(Z2F,cccccccccc
cc	ccc
	c
	cP(V<VF(<P(((F(P222Z<PP2FZ2(<<<Z(<P2F<<<	cc
c	ccccc	c	c
cc5		423454234235544446798987BX*\$b<X"\(`�<BZ(R$X<Z"`x,R<"Z�$\NV ^(P2Z,TFdNnLl,TDvNd<X(FZ<^ * *^	cc
cc	cc
ccccccc	%%%%&&&&''''%&%&P(<ZDP<
Z$2(."rfnd
($""""RDbPb"h$2P
Vcc	ccccccccccccc	cccccc	c	cc
cc(	 #!"( #%&%&%&( "#( "#!F`6(0\D$$P"F(Z<
PF&"<8P: 2Z(PZjf"`Z<P
Z <P"Z(<<"$"Z<P(&%(Z<(222(<Z(P(P2<(Z2 ��	
  ����  ��  ��������(((&*.$(8HXh @������߿	   	 	$-5;?BDGHGDB?;5-$	 ,BXn������6Lbx �� � � � � ����� �Ԙؘ֘ژܘޘ����������� �&�,�2�'!))+1	-9
/=		
12354

��   �    �
$%<<<<<<<<<<< ���  ��   �����Ιљԙי��ϙә֙ޙ��Йҙՙ����c'(c
'c`'*+*+-.c' ' ' >>>>>>c((c''(P 

	






           	
& #678999	
@

	9A ����}2�dd�PP8 3<=> :;CDEFGH22d������





 "$&����������  ��  ����  0@P`p��������  0@P`p��������  0@P`p������������������������������������������? �� ��� �    �? ���?     �?<  �   0�  ����  0      � �  �?� ��     0   ���>ë����������? ��������:  �  �� �   �  ��   ������������������������������������   �    � �      � ������������������������������    �����   ��   �  �     ������������     � �����������    � ����������������    �     ��������  � ������ � ������� �    �  �    � � �� � ������< ����  �0   �?  0 ?  �����������0 �*�0 �� * �  ����� �� � � �� �������ꯪ��   �  �    �   ª����ꪪ��   ����   0�����?�� �� ���  0     0   ����  ��    ��   �����  � �  �     �꺪�  �  8���  ȃ ê�������0� �<� ������� ȃ�������ꪪ�� (� �����������V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V���        7�� �p3� L��U\uU�zU� ������ �?        ��:�  <   �  ��  0 � ����Uu<�Zu0L<�Zu�Uu ��� 0 � ��   �   <       <   �  ��  0 � ����Uu<�Zu0L<�Zu�Uu ��� 0 � ��   �   <                     � �������� ��?                             � ? � <� 0< <� 0�<� ��������?�?<��� �?  0�  <�� �    ?�?  �  < ���?  �����3�?3�? ��?� ���?<�� �0�< �������0�? �� �  < ���?  �����3�?3�? ��?� ���?<����0� �� ��?  ��  �� <?  ��?���0���0���0 �����?�?��<���0������ ����?�0<     �  < �< 0<0 <0  � <����  ��?0< �?<�?0��  �?� ? �? p� \��_�����_|]�� �?    <<���<<     ��         �  �< ��� �����?<<3����:� 0�� ��  ̨ 0� ��6 �� 0� ��   �  �  p�  _� ��� � ?� ���*� �� � ? ���  _�  p�  �  �       �   � ? ����:�����UU��������������
��
������������������������������������������������                    <�                    ��                    <��������������������������?�?����������VU�VU�������
*������VU�VU�VY�Vj�������������VU�VU��U�������������0 ���VU�VU��i��i�������������VU�VU�������
*�����V�Z�h)�
������ �U�hii
ZZZ)��V)hUU
�U��U� ��� �U� �U� ��� �U�h�Z
ZUU)���*  � �   �  0  �?  0 �   � �� �3 �? ?� \��� �W0�  0� �s0���  p��/ p�?��  p�� 02 𨪪  Q03  �Q�    0  ����:   2�+0   ��+�  �?��/�  ��0 ?�  <�� �0  < � �0  � � ��  � ��  �< ��   <  <    < (3    < (3    ? (3    ? (?  (�(�*���

(�(
�
� � �
�
�(�(��

�*�     �? �� ��<�,���:��? �� ��  ��  �      <   0   0������������UUUUUUUUUUUU��������������������������������������������UUUUUUUUUUUUUUUU��������������������������������������������������������UUUUUUUUUUUUUUUUUUUU  �?    �?    �?    �    �?    �?    �?   ���   ���   �?�   �?�  ��  ��  ��  ��  ���  ���?  ���?  � �? �� �� �?  � �?  � �?  ��� ��?�� ��?�� ��?��   ��   ��   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �?   ����� ���? ��� ����������? �? �? �? �? �? �? �? �? �? �? �? �? �? �? �? �? �? �? �? �������  ��  ��  �� �� ��? ��? ��� ��� ���������������?�� ?�� ��� ��� ��� 0�� ���  ��  ��  ��  ��  ��  � ����������������  �   �   �   �   �   �   �������������   �   �   �   �   �   �   �  ������������ ���0 �?3�3 3��?0   0<����<�0   0 �<����0<           00     <0�   �   � �   0�*�   � �  ����   < �?<    �?�  ���  �?���  0��   <�
��  ̬
�:   ���
? �?��*�   ����   �����   � ���  0 � �   , � 0   ,� �?  ���  ��|�  0?�@�  �?P�   �@� � �5� ��1�?� |u�� ��V�����VUUU�VUUU�VUUU�VUUU�VUUU�VUUU��������V�V�V�V�V�V�V�V�V�V�V�V�V�V�����j�Z�h)h)�
�����
h)h)Z�j��� 
( �*� ���h�V
ZiZ)�������jZUUiZUUiZUUiZUUi���j����ZiZ)h�V
����*�  
(      �        L% �]I �qH@f6 P* ��� P ,j��#@$�(  ��f  �Z ��f       0     �      ��    �      0    �      �� �   �?  ���*VU 3 
��
 ���/   ���:  �
��    ����     ���     ��:     ��      �      �(      ��       
           �     �
     ��      �+      �*      �     ��     ��     *�    ����    ����             ���    ���*  �����*  �����* ������?  �  �:   X����� �V����� hը���� X5�   �گ��*�`=������+���*��*��   �*�����:������� �� ��  ꪪ�� ��
  � �ꪪ��  ꪪ��
  �    �    �   �0� �0  �?  � � ?  �  �3 �� 
?�  ?<  �� �? ������               �                            �   � < à    ����     �*
   �#�   �$�   �P%��	  <h� D+  ��	 "  8   ���
���           ��(  ��( hiW  *Z  �  ��  E�   ��� I*   �/@�
   �<& 
    ����+   �+0!�/�   
�+   � �
+  (���    
8�
�    � 0       <        2    �? �  ���  ?�0 ��� < ��
� �   ��  * �� �* �����
 ��(�( �*�"
ª����
������������������ ?        �����   ?   ?�<�� �3  �� <�+< ��   �*��?��    �� � �     ��? � ��  ��  � � �  ��.�?  � �  �    � �* ���   �� �*
  �� ��� ��* ��ꫫ
 �� ��?�����  ����������
 < ����������
������������� �����������������������������������   �  ��? �� ��Ϫ��>���;���;����������>������ �������
��
 **  �
� ��� �� ����������������  <  <0 �  �� �  ���� ���� ���� ���� .��� +�����+�����*�����*�����*�ϯ��
������+�� +��< ���
��� � �*����
�/���*ꪪ��
������������ �?   ��   �&  � ��* Ͼ� ÿ" �*> ��< �
< �*< 
���  �� �� �� �
�  ��� �����*��
 � �� �� � ;  � ?  *  #
  "*  "
  "
   �      �
   ��� �*
(��* (�� ��*��
�������������  *    �  �*  U� �WU��pUU)�_UUT� ���������*����  ��� 
�����*�� �
*
������ ��������������������������    0 ��  �?  0<�0�������� <<3��?����� ���?̺*������
�*���
�� �� �
�*���      < 0 � � ?  <3  <  ?�? <� � 30���3� ����0� ��?� ? ��<����� �
"  �� ��
�*
� ������*�  ����
�(
���������   �0 �(���0
������?��������������
�?*�<:�����(����*������� <��
<������� �+�0 ����2�
���
��������*�����             � 0    0  0 �   0 ��   < ��?  � ���< ? � � ��� 0��������3�< * ���0����?�� ����� �? 0�( �  � ��� �  � ����>� �*�
���(2 ��
�
*�����(
������������������ 0     ?  ��? ����  <��  ���<<��*�� ��� ��+���+0����0� ���? ����   �0  ��*0�  ���?  ���0 � ��������((�����"������  � �   ��  � �� ( <�� ( �?0* ��  3���? ��� ��� / � �+�3 ���� ������( "�����(��(*�
������H�� �P�� ݩ$�� �� �� �� �d�� ݩ� �q�� ݩ� �~�� �h`H�� �d��v  bܭu  bܭt  bܩ� �q��y  bܭx  bܭw  bܩ� �~��|  bܭ{  bܭz  b�h`H�Z�q �| �N��p �{ �D��o �z �:�q �y �P��p �x �F��o �w �<�q �v �J��p �u �@��o �t �6��I ε � ��b� �} ������� �- 4��b� �� ������� � ε !��b� �� ������� z�h`�w �z �x �{ �y �| � �� �� ����`�t �w �u �x �v �y � �} �� ����`�o �t �p �u �q �v `�o �w �p �x �q �y `�o �z �p �{ �q �| `H�Z�� � �L� �� ϴ����� �b�% ���%H�a�%���  }� ��h�%���  }ܭ  ��������%�b� g�L϶�
�%L϶����%�b� ��L϶�#�%L϶�� B��C B�Lh���� ����  }�� ��� �Lh����Lh� ����  }������ �Lh��� z�h`Z�� ��
��	�� ȹ	�� ����b�8�7��b�%z`Z�
��	�� ȹ	�� ���%�b�i7��b�z`H�Z8�7��%�a�
��%��A8�7�%��a�%h`H�A8�7��%�a���0�%��Z8�7�%��a�%h`H�����h`Hڜt �u �v �w �x �y �z �{ �| � �b�} �� �� ����$�} �� �� �h`} � � dq~                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���ة��  ��� � �� � �� �ߍ& ��" � t ���� �� �� � ����� ��� ��XL �H�Z�����������������
��
�	��	���������������� ��������� �a��a���� ���ރ����� ��� � :� �z�(h@H�' )���# �$ �% (hX@                                                                                                                                                                                                                                          �휏 ���$���&   ��ߍ& � K񩖍�  ����� ̷ �� C� �� ?� ���`��<�l�o �p �q �r �s � �b�u��^�]�s�t��n�o�m�,�+�h�i�j�k�>�?�V �:�=�;�*�v�* �+ ���# �@�) ������	�
������' ��� �4�0�d�k�" �	 � ���������$���a�)��q�+�\� �$ ��% �� � �$����% ����_�'` �� �� �� ������'����' �ĭ��� C� �� C� �� �� �� �� �� M� ǩ  �� +ĭ��  ��a �� �� ��� �ƭl��J���  ������7�t���0������з���<� }� �ĭ`�H���< �� �ƀ� ?耐` |�`���m�� �� � �� � #� �ʩ� ��`�� �� -� �Ω� K� � T� ͌ � �� ��`��6 �� �߭t���� � ,� m� Ԇ �� � ���  �� Q٩�`H C©�l vÜlh` ��H�` �� Eũ ǭ  ��`����u������u �� � cŭu���V��H�` Eŀȩ� ��� �ڢʽt  b�� ���� ��� ݢʽo  b�� ����� �F�� ݩ� �T�� �`�
� �`���!��"��  L�`�
� �`���!��" C�` ��� �(�� ݩ� �<�� ݩ �`H�
� �F��l��i
 ݩ�"�X�# |ǩ �h`Hڭt����&���:��o mr �o �p ms �p �q i �q ؜r �s �� ����ʽo  b�� ���h`H�Z �� �� �� ��  ���)��&  �� �Ʃ� ����	 ݮ  ��� �� �� �� �� �� ��ߍ&  �� 7���� �� �  K�z�h`H� � ����(�!��" C�h`�t����	��]�]�F����&���	`�&���� � ���l�l�� �Ɯ&`� �ũ � ��&��� K Z� �� ���"�P�# |ǩ  ��` �� ������`H�l��F��"�P�# |ǩ � �̭"���"�� |ǩ ǭ"�� ���"��%�e�f�gh`��"�P�# |� t�h`H��!��"�� �"� �#� L�h` �� ��`�l���  ���X��� ƀO�� �̉� �̉� �̉� �̉ � ȀH�;� !� �� wȜ;h�� ȀH�' ����' h�@`H�' h`H�;�;�0 ��h`H ��;�0
 � K�h` ��h`HZ� �,� �4����g  ���g zh`HZ� �D� �L����g  ���g zh`H�m�� ��h`H�"� =�* �8�+ �3�- �"i��#i� gɜ, �"i��#i� �� ��h`Hڭ* �� �`�,* � *����� ;��h`Hڭ* �� �`�,* � K������h`Hڭ* ��* �9�- � �,��4� g��h`H�,� �4���!��"��  L�h`H�,� �4���!��" C�h`Hڢ �- ���. �ɭ- ���$��,��4�`�* �* � ��- �9�����h`�- � �ɀ�� ʀ�� Mʀ�� ��`Z�iɐ����  B� A��
� U���z`���- z`��-  ��z`Z�i�':� �� B� A��
�� A��
�� �z`��-  ��z`� ��- z`���- z`Z8��05���  B� A�ȱ$�
���z`��-  ��z`����- z`���- z`Z8��0F� �� B� A��$�
�� A��$�
�� �z`��-  M�z`� ���- z`���- z`Hڭ+ �� �`�,+ � G����� Y��h`Hڭ+ �� �`�,+ � h������h`Hڭ+ ��+ �8�, � �D��L� ���h`H�D� �L���!��"��  L�h`H�D� �L���!��" C�h`Hڢ  �˭, ���$��D��L�`�+ �+ � ��, �8�����h`�, � �ˀ�� ̀�� Q�`Z8��0���  B� A��
� U���z`���, z`��,  ��z`Z�i�'� �� B� A��
�� A��
�� �z`��,  ��z`� ��, z`Z�iɐ�+���  B�� A��
���z`����, z`���, z`H��f�ih`H��e�hh`H��j�gh`H��%�+h`H �� � |� ����� Y�h`H��!��"�"� �#� C�h`�% I͜%�e I͜e�f I͜f�g I͜g`�l�� {� �̭,���# ���"i�(�#i�)���g  ���g  J�`Z��_�m"���"0�"���"�d�m#�#�#����#z`H��0�a��� �̭#���a�_� �̭#�l����a�_��h`�"� � �#i� B� ����D� ����:�l���i��"� ��#i��"� �  B� ����� �`�Z A��9�
�1�1-���� ���
� �� ���m� t��m�m����m����� z�`H�_�% �̩�"�?�  Lݩ *� � Cީ����_h`HڭV ���;�"�"/� �`�,V ����%��V �V �"i�W �#i�_  � ���  *��h`HڭV �&� �`�,V � ������`�,V � �������h`HڭV �&� �`�,V � a������`�,V � �������h`HڭV �� �`�,V � J������h`HZ���
�>���'�4� ������9��!�h��"����  Lݭ�! h� ����� Y�zh` ��zh`HZ���(� ������9��!�h��" �� C�zh`HZފ04������������� йB�}���������
� ��� ��zh`�������u �`H�! ���'�� cН�� ��h`Hފ0)��������� cН������� Щ ��� ��h`��� ��� B� A��
����� U���`HZ��0#���� й.�}���8��� �������������zh`HZ _����iJ�� � A��
����� U�����j� ���! �� �zh`H��!��"�� �i� �j� Lݩ��kh`H��!��"�i� �j� Cޜkh`HZ��� �����!��"��  h� Lݭk��� +�zh`HZ��i�x�
��� /Ѐ
���<0 �zh`HZ8���0�����@�}������ ��zh`H�
��� �����h`Hފ ��h`HZ��� �����!��"�m�䐍  L��! h� ��zh`���4� ��`� ��`H������ފ�3�� �Ҝ+�� �����+�(� ���2�� ����� �Ҝ+h`H�����<����(����
���� ��h`HZ��i������^��ҍu ��^�^���^zh`H������ފ��� �Ҝ+��Ȱ �Ҁ�
��h`������ z��! 
��� ȹ� � �}�� ����}�� �� ��`HZފ0���������zh` ��zh`HZ�! �� _����iJ�� � A��
����� U�����j� �� �zh`HZ���
��i���:�06������ z��! 
��� ȹ� � �}�����}��������<� ��zh`HZ��
���$ ȹ�% � �$}�� �.�(�*����$}������ �ɀ����������zh` ��zh`HZ���"���� ��� �����������zh`HZ���"���� ��� �����������zh`HZ���"0���� ��� �����������zh`H��ɂ�� �� �Խ���&��h`H����ފ�1����
�����#�8�����������i�l��l���������+��<��+��n��+���������,� �Ҁ ҂h`HZ8�����\�}�� ��'����`�}�� �	ɀ���� ��zh`H�����
T��iɐ1��h`H�����
:ފ0h`H�����
(8���� ���� ��h`H�����
	���'������� z��! ���$��h`HZ��
���$ ȹ�% � �$}�0�'����$}�� �
�n���zh` ��zh`H�����(� ���)�
0 ���iɐ�靜�8�����ڝ�ފ0�h`H�����(� ���)�
0 �8�����靜���iɐ�ڝ�ފ0�h`H�����
���i���ފ ��h`H���*ފ������L����i�x����L�ם�L����)ފ��������m8����
�� ��L�ם�L����(�����$�� ��L����i�x�����.���)��%�����$�����8�����������h`H�����ފL��8�����L��"ފL��$8�����L��?��i��L��Lފ�/�g8������ �l����{��i���ފ ��h`H�������L���8�����L�����L���8�����L���9��i��L���H���4�b8������%�gފ��w��i��������'0 ��h`H�Z����� �`�,������� ��z�h`HZ�! ��6�8�2������'�� _���� �zh` kڜ\zh`Hڭ�� �`�,� ������h`Hڭ�0� �`�,�
��6�
 <������2�\�\�80���\��h`Hڭ�/�\��� ۢ �`�,�
�i2�( ������ ����� Y��h`H�Z��� � ���6�� ���h�-��>�':���8��2�����!���"��� ��50�
�( =� �٭�! h�z�h`� �4� ��` ��`HZ���(+� � � ���8��2�����!���"�! C� ��zh`HZ����5� �7���������u ��2�zh`H�&�2��3� �6��7�5��� ��h`H�Z�7�� �6 ��� ���i������ ����6��z�h`
m5����p�m2������P���!8� ������m3����6��u �`H�5�5���5�6�6���6�7�7���7 ��h`H� 
��F�� ȹF�� �!�#��"� � � 0m!�)008�(� �#��"8�!�m � � i � ��#�� ���m � ���i � h`HZ� �!�� ;�� � i � ��#�#�#8������4�NnNn����ȱ���� ��!���  ���zh`�4� ��` ��`H���4���NN����h`Hڪ)�JJJJ�% }܊)�% }��h`xH�Z�%�a��$��b��%��c��&��d��'��d�� ���� ��#���� ���� � �-$�� i� � i � Ȳ-$�� i� � i � ��#к� � z�hX`H�Z
��+��$ �+��% � �$�$�&�a��b��Z0��b��0�b�8�7�% }�Ȁ�z�h`H�Z� 
��F�� �F�� �!�#��"� � � 0m!�)2�l�� 06�`�!m �#�8� � � � � � � � �<8�(� �#��.� m� � m!� � i � ���8���� � ���m � ���i � � ����#��� m!� � i � � i0� � i � � ��� ��z�h`H�Z�!�#�"� � � 0m!�(�;�� 0�/�!m �#� � � 8�(� �#�� m� 8���� � ���m � ���i � � � ���#��� i0� � i � � ��z�h`H�Z�  	����� � �� 	߭t��� �� ����� Y�z�h`Z�. �!�6 �"�> � �F ��N �$��  �� ��l�0� ����c �� ���cz`H�Z� �. �!�6 �"�> � �F ��N �$��  �� �߭l�0� ����c �� �ߜc� �	��е� ��z�h`H�Z� �. �!�6 �"�> � �F � �� S�l�0� � ���  S�� �	���â ��z�h`HZ� �#�	��Ȁ�� � ���zh`HZ� m!� � i � �c���� i0� � i � zh`8� �0� � � � zh`HZ�#�#� �#� �Ȁ�� �� i0� � i � ��zh`HZ� 
��F�� ȹF�� �!�#�"� � �8�!�
 m � � i � �
 �#�� �
8�!� �#�c���
�m"�����m � ���i � zh`H� � �߀ M�h`H��� ���NN����h`� � i � �
 �#�#`HZ� � � � 7��#8������ �NnNn����ȱ���� �� ��  ���zh`Hڮ �. ��6 �� � � � � � � � � ���N.N.������&� m� � i � � i0� � i � L���h`Hڮ �. ��6 �� � � � � � � � ����NnNn������&� m� � i � � i0� � i � LQ��h`H ��l�0 (� �� � i � h`H�t���� ��
 � e�� � �� ��� Ԇ ��h`H�Z�>� �	 � � � �l
��� ȹ� � ���N�	 �> � ��. y> �	 ���6 8���6 �F �	 �*	� � Ȁɮ �. �
 � �. �  �z�h`Hڮ �. �!�6 �"�> � �F � ��� � ��� � �. �
 � �h`H�Z� �l
��� ȹ� � ���c�� �" �n�o���t� ���2� � ��� � �N� ��. � ���6 8���6 �F �(�>  �z�h`H�Z� �F ��i'� ���i � � ��i'� ���i � �N �$�
��F�� ȹF�� z�h`H�
 � e�� � �� M�h`Hڮ � �> ���� �> � ����h`H��  �����
0�h`H�  ����h`Z����z`Pd������Z�� �� ���z�`H�Z� �@� � � � ����� ���� �z�h`H�� 3���
� +�<�
�� ����� I�
�h`Hڭ���� �`�,������	��� Q��h`H�" ��������� ������ ��������" �" ���" h`Hڭ��"� �`�,�� �� ��`�,�� �������h`HZ��� ������8��!�>��" C�zh`HZ��� ������8��!�>��"�D��  L�zh`H�����i����(������ފ��h`�h�-���h`H 5������ ��h`HZ�u���Q�!�J��!��"�O�� �T�� �X� L݀�8���Y�� �[���]� ��u�u�zh`���uzh`�  ���]�]� ����'zh`����'zh`H�� ������h`HZ�
����$ ȹ��% � ��!�$� ȱ$�"ȱ$� ȱ$� L�ȱ$�  L�� ��"ȱ$�!��$�  L�zh`HZ��H
����$ ȹ��% ��$�"ȱ$� ȱ$���! C�ȱ$�  Cީ�"ȱ$�!��$�  C�zh`Hک � ���� ݩ � ���� ݩ� ����ʽo  b�� ���� � ݩ� �����!��"��  Lݜ��<� ������h`HZ��.�� �����!��"��  L�zh`HZ�<�.�� �����!��" C�zh`H�  �� ��� �P�� ݩ � Z� �� �� M��< ���"�P�# |�h`H�l��4 �� �� &��
� �� � ��P��7�� � G��� � �� �h`HZ�=��#�=i� �����!��"��  L��=zh`H��!�� �����" Cޜ=h`H�0 ��h`�W �'� �_ ���!��" ���& ����h�-V �V h`��  L�h`H�W �W �'0	�h�-V �V h`H�0 ��h`�W � �_ ���!��" C�h`H�W �'-� �_ ���!��"���g  ���g �& ���
�=�  L�h`�h�-V �V h`H�W � �_ ���!��" C�h`Hڭ)���&��`�,V ������V �V �(i�W �)�_ �h`Hڢ�`�,V ������V �V �"i�W �#�_ �h`�
�����$ ȹ���% ��$`�(� �)����g  ���g �& `H�\�)� �( J쩪�,h`H���)��� �� �� Y� J�
�h`�,ɪ��(i�(�0R�,�M�' ���+�,��� M�q���
 6�s���+ ��& ���' �,��,����q���
 6�s��� �`�+ 5�+�h 5�h�i 5�i�j 5�j`Z��_�m(�(�d�m)�)z`HZ ���(��)� z��! 
��� ȹ� � �m(�(��m)�) Y���� � J�zh`�"�(Fi�(`8�#�)0��)0`�#i�)` ���"i�(8�#��) J�' ���,`8�"����(0`8�#�)0��)0`�#i�)` ��8�"��(8�#��) J�' ���,`Hh``8`` ��`8`8`` ��`HZ�(� �(�	�'0�'�(� �)� ���)�	ɀ����)���!��"�*�%��  L��*�*���*zh`H�Z� ��l ��#��k � ���� ���� �k �-$�l ��k �k �(�� i(� � i � �k ���m ��l �Ŝ� �l ���n Ф�� �#�z�h`Hڍ� �� ���� �h`H�Z�� ���F�� 
����� 轕�� �� 

����'�* ȱ�



�� �� ȱȍ� �) ȱ�� �( �� � ��z�h`�� �* `������    
 (	� # � �� ��  �� �� � � � � � � � �� �� �� �� �* �� �� �ߍ& `H�Z�� ���Q�� ���.�� � �� �� � �  �ﭭ � �� �� � �  7�� �� ͛ � ��� �� ͨ � uﭕ ���.�� � �� �� �� � � � �  ��� �� ͵ � �z�h`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
����� ���� Ȍ� �� �� �� � �'�� ���� ȱ��� � ��� � ��� ��Ȍ� �� ��`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
����� ���� Ȍ� �� �� �� � �#� ��  �� �� �� � � �� �� � � `�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
����� ���� Ȍ� �� �� �� � �'�� ���� ȱ��� � ��� � ��� ��Ȍ� �� ��`H�Z�� )?	@�� �� 4��-� �� �� ����� )@��J��� �� Ȍ� �����Ρ �� �� �� Ϳ �� �� z�h`H�Z�� )?	@�� �� 4��-� �� �� ����� )@��J��� �� Ȍ� �����ή �� �� �� �� �� �� z�h`H�Z�� )?	@�� �� 4��-� �� �� ����� )@��J��� �� Ȍ� �����λ �� �� �� � � �� �� z�h`� �� `� �� `

������ ȹ���� ȹ���� ȹ���� � ���� ���� ȱ��� ���� �� �� ��� ��  �� u� �� 7���� `�ZH
������ ȹ���� �� ���  � ����� hz�` �  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  w�     q�  j�  d�  K�  Y�  K�  Y�  w�  ��  ��  �� .� }� }� �  ��  ��  j�  Y�     q�  ��  ��  ��  ��  ��  ��  �  _�  K�  ��  d�  _�  T�  q�  d�  _�  q�  �  ��  ��  ��  ��  ��  �  ��  �     �  q�  d�  q�  ��  ��  T�  _�  T�  K�  _�  ?�  G�  G�  T�  G�  d�  T�  _�     ��� ���.���.��.�@�.�@�h�@�@�T�� ��� �� �� �� ��    _�  Y�  T�  O�  K�  G�  C�  ?�  ;�  8�  5�  2�  %�  ,�  ;�  K�  _�  w�  ��  ��  ��  ��  j�  O�    ��T� ��T���T� ��T���T� ��T���T� ��T�T� �� �� ��T� �� �� ��T� �� �� ��T� �� �� ��   }� �� �� ��}� �� �� �� ��T� ��T� ��T� ��T���T� ��T�T���   T���T���T���T���T���T���T���T� �� �� ��   ����������������������������������������������������������������   ��������������������������������������������   ������������������������������������    *� /� 8� ?� T� _� q� � �� �� �� ��T�}�����   ������\�����}�T�.� �� �� �� �� �� � q� _� T� K� ?� 8� /� *� %�    *� /� 8� ?�T� _� q� �    *� /� 8� ?� T� _� q� � �� �� �� ��T�}�����   ������\�����}�T�.� �� �� �� �� �� � q� _� T� K� ?� 8� /� *�    ��.� �.� �� ��.� � �� �
� �
� �
�T� �}�T�.�� �T�.� �
�.
� �
� �
� �
� �
� �
� �
� �
� ��    � �� �� _� T� �� � �
� �
� �
� ��   ��\�\�\�\�\�\�����\�\�\�\�\����
��
��
���������\�\�\�\�����\�\�\�\�\�   \���\��
�\
��
��
��
��
��
��
��
�\�\�\�\���\�\�\�\�\�\�}�T�\� ����
�\
��
���	    U�   h�������������������:��\��������������     �� /2�	    �

� �	
	 �				� �	��				 �

		����������������������������$�  ��$���  t���.��  ��      ��E�  ��  ��>�  ��>�  ��R�  ��4�  ����#�$�  1�7�B�J�Q�^�c�l�q�w� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____xH�Z�h 
���� ��i@� �m �#�n ����� ���� � JJ��-$�� i� � i � ��� �Ȁ��#�#� �
�n ��L��z�hX`H� �$ m����$h`H�Z�/���� ���� ��z�h`�`�a                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           O� ���